`ifndef ASIC_DEFINES_VH
`define ASIC_DEFINES_VH

`define XLEN 64
`define EXTMEM_ADDR_SIZE 24

`endif
